Unid