-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.0.0 Build 614 04/24/2018 SJ Lite Edition
-- Created on Mon Sep 24 17:34:28 2018

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SM1 IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        Z : IN STD_LOGIC := '0';
        proximo : IN STD_LOGIC := '0';
        enable : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
        selectTempo : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        selectConstante : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        selectFuncaoULA : OUT STD_LOGIC;
        resetReg : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
    );
END SM1;

ARCHITECTURE BEHAVIOR OF SM1 IS
    TYPE type_fstate IS (cus,mais_us,cds,mais_ds,cum,mais_um,cdm,mais_dm,cdh_2,cuh_4,cuh_9,mais_uh,mais_dh,nada);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,Z,proximo)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= cus;
            enable <= "000000";
            selectTempo <= "000";
            selectConstante <= "000";
            selectFuncaoULA <= '0';
            resetReg <= "000000";
        ELSE
            enable <= "000000";
            selectTempo <= "000";
            selectConstante <= "000";
            selectFuncaoULA <= '0';
            resetReg <= "000000";
            CASE fstate IS
                WHEN cus =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= mais_us;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= cds;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cus;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "000";

                    selectFuncaoULA <= '1';

                    selectConstante <= "100";

                    resetReg <= "000001";
                WHEN mais_us =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_us;
                    END IF;

                    enable <= "000001";

                    selectTempo <= "000";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN cds =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= mais_ds;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= cum;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cds;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "001";

                    selectFuncaoULA <= '1';

                    selectConstante <= "011";

                    resetReg <= "000010";
                WHEN mais_ds =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_ds;
                    END IF;

                    enable <= "000010";

                    selectTempo <= "001";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN cum =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= mais_um;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= cdm;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cum;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "010";

                    selectFuncaoULA <= '1';

                    selectConstante <= "100";

                    resetReg <= "000100";
                WHEN mais_um =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_um;
                    END IF;

                    enable <= "000100";

                    selectTempo <= "010";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN cdm =>
                    IF ((Z = '1')) THEN
                        reg_fstate <= cdh_2;
                    ELSIF ((Z = '0')) THEN
                        reg_fstate <= mais_dm;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cdm;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "011";

                    selectFuncaoULA <= '1';

                    selectConstante <= "011";

                    resetReg <= "001000";
                WHEN mais_dm =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_dm;
                    END IF;

                    enable <= "001000";

                    selectTempo <= "011";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN cdh_2 =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= cuh_9;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= cuh_4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cdh_2;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "101";

                    selectFuncaoULA <= '1';

                    selectConstante <= "001";

                    resetReg <= "000000";
                WHEN cuh_4 =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= mais_uh;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cuh_4;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "100";

                    selectFuncaoULA <= '1';

                    selectConstante <= "010";

                    resetReg <= "110000";
                WHEN cuh_9 =>
                    IF ((Z = '0')) THEN
                        reg_fstate <= mais_uh;
                    ELSIF ((Z = '1')) THEN
                        reg_fstate <= mais_dh;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= cuh_9;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "100";

                    selectFuncaoULA <= '1';

                    selectConstante <= "100";

                    resetReg <= "010000";
                WHEN mais_uh =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_uh;
                    END IF;

                    enable <= "010000";

                    selectTempo <= "100";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN mais_dh =>
                    IF ((proximo = '0')) THEN
                        reg_fstate <= nada;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= mais_dh;
                    END IF;

                    enable <= "100000";

                    selectTempo <= "101";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN nada =>
                    IF ((proximo = '1')) THEN
                        reg_fstate <= cus;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= nada;
                    END IF;

                    enable <= "000000";

                    selectTempo <= "000";

                    selectFuncaoULA <= '0';

                    selectConstante <= "000";

                    resetReg <= "000000";
                WHEN OTHERS => 
                    enable <= "XXXXXX";
                    selectTempo <= "XXX";
                    selectConstante <= "XXX";
                    selectFuncaoULA <= 'X';
                    resetReg <= "XXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;